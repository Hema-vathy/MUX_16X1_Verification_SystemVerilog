//files block
package file_pkg;
`include "clock.sv"
`include "reset.sv"
`include "stimuli.sv"
`include "rst_test.sv"
`include "comparison_test.sv"
`include "run_test.sv"
endpackage
